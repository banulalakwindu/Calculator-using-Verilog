module Divider(input A6,A5,A4,A3,A2,A1,A0,B6,B5,B4,B3,B2,B1,B0, output Q6,Q5,Q4,Q3,Q2,Q1,Q0);

UnitCell u1(A6,B0,1'b0,u2_sout,u1_out,u1_bout,u1_sout);
UnitCell u2(1'b0,B1,u1_bout,u3_sout,u2_out,u2_bout,u2_sout);
UnitCell u3(1'b0,B2,u2_bout,u4_sout,u3_out,u3_bout,u3_sout);
UnitCell u4(1'b0,B3,u3_bout,u5_sout,u4_out,u4_bout,u4_sout);
UnitCell u5(1'b0,B4,u4_bout,u6_sout,u5_out,u5_bout,u5_sout);
UnitCell u6(1'b0,B5,u5_bout,u7_sout,u6_out,u6_bout,u6_sout);
UnitCell u7(1'b0,B6,u6_bout,~u7_bout,u7_out,u7_bout,u7_sout);

assign Q6 = ~u7_bout;

UnitCell u8(A5,B0,1'b0,u9_sout,u8_out,u8_bout,u8_sout);
UnitCell u9(u1_out,B1,u8_bout,u10_sout,u9_out,u9_bout,u9_sout);
UnitCell u10(u2_out,B2,u9_bout,u11_sout,u10_out,u10_bout,u10_sout);
UnitCell u11(u3_out,B3,u10_bout,u12_sout,u11_out,u11_bout,u11_sout);
UnitCell u12(u4_out,B4,u11_bout,u13_sout,u12_out,u12_bout,u12_sout);
UnitCell u13(u5_out,B5,u12_bout,u14_sout,u13_out,u13_bout,u13_sout);
UnitCell u14(u6_out,B6,u13_bout,u15_sout,u14_out,u14_bout,u14_sout);
UnitCell u15(u7_out,1'b0,u14_bout,~u15_bout,u15_out,u15_bout,u15_sout);

assign Q5 = ~u15_bout;

UnitCell u16(A4,B0,1'b0,u17_sout,u16_out,u16_bout,u16_sout);
UnitCell u17(u8_out,B1,u16_bout,u18_sout,u17_out,u17_bout,u17_sout);
UnitCell u18(u9_out,B2,u17_bout,u19_sout,u18_out,u18_bout,u18_sout);
UnitCell u19(u10_out,B3,u18_bout,u20_sout,u19_out,u19_bout,u19_sout);
UnitCell u20(u11_out,B4,u19_bout,u21_sout,u20_out,u20_bout,u20_sout);
UnitCell u21(u12_out,B5,u20_bout,u22_sout,u21_out,u21_bout,u21_sout);
UnitCell u22(u13_out,B6,u21_bout,u23_sout,u22_out,u22_bout,u22_sout);
UnitCell u23(u14_out,1'b0,u22_bout,~u23_bout,u23_out,u23_bout,u23_sout);

assign Q4 = ~u23_bout;

UnitCell u24(A3,B0,1'b0,u25_sout,u24_out,u24_bout,u24_sout);
UnitCell u25(u16_out,B1,u24_bout,u26_sout,u25_out,u25_bout,u25_sout);
UnitCell u26(u17_out,B2,u25_bout,u27_sout,u26_out,u26_bout,u26_sout);
UnitCell u27(u18_out,B3,u26_bout,u28_sout,u27_out,u27_bout,u27_sout);
UnitCell u28(u19_out,B4,u27_bout,u29_sout,u28_out,u28_bout,u28_sout);
UnitCell u29(u20_out,B5,u28_bout,u30_sout,u29_out,u29_bout,u29_sout);
UnitCell u30(u21_out,B6,u29_bout,u31_sout,u30_out,u30_bout,u30_sout);
UnitCell u31(u22_out,1'b0,u30_bout,~u31_bout,u31_out,u31_bout,u31_sout);

assign Q3 = ~u31_bout;

UnitCell u32(A2,B0,1'b0,u33_sout,u32_out,u32_bout,u32_sout);
UnitCell u33(u24_out,B1,u32_bout,u34_sout,u33_out,u33_bout,u33_sout);
UnitCell u34(u25_out,B2,u33_bout,u35_sout,u34_out,u34_bout,u34_sout);
UnitCell u35(u26_out,B3,u34_bout,u36_sout,u35_out,u35_bout,u35_sout);
UnitCell u36(u27_out,B4,u35_bout,u37_sout,u36_out,u36_bout,u36_sout);
UnitCell u37(u28_out,B5,u36_bout,u38_sout,u37_out,u37_bout,u37_sout);
UnitCell u38(u29_out,B6,u37_bout,u39_sout,u38_out,u38_bout,u38_sout);
UnitCell u39(u30_out,1'b0,u38_bout,~u39_bout,u39_out,u39_bout,u39_sout);

assign Q2 = ~u39_bout;

UnitCell u40(A1,B0,1'b0,u41_sout,u40_out,u40_bout,u40_sout);
UnitCell u41(u32_out,B1,u40_bout,u42_sout,u41_out,u41_bout,u41_sout);
UnitCell u42(u33_out,B2,u41_bout,u43_sout,u42_out,u42_bout,u42_sout);
UnitCell u43(u34_out,B3,u42_bout,u44_sout,u43_out,u43_bout,u43_sout);
UnitCell u44(u35_out,B4,u43_bout,u45_sout,u44_out,u44_bout,u44_sout);
UnitCell u45(u36_out,B5,u44_bout,u46_sout,u45_out,u45_bout,u45_sout);
UnitCell u46(u37_out,B6,u45_bout,u47_sout,u46_out,u46_bout,u46_sout);
UnitCell u47(u38_out,1'b0,u46_bout,~u47_bout,u47_out,u47_bout,u47_sout);

assign Q1 = ~u47_bout;

UnitCell u48(A0,B0,1'b0,u49_sout,u48_out,u48_bout,u48_sout);
UnitCell u49(u40_out,B1,u48_bout,u50_sout,u49_out,u49_bout,u49_sout);
UnitCell u50(u41_out,B2,u49_bout,u51_sout,u50_out,u50_bout,u50_sout);
UnitCell u51(u42_out,B3,u50_bout,u52_sout,u51_out,u51_bout,u51_sout);
UnitCell u52(u43_out,B4,u51_bout,u53_sout,u52_out,u52_bout,u52_sout);
UnitCell u53(u44_out,B5,u52_bout,u54_sout,u53_out,u53_bout,u53_sout);
UnitCell u54(u45_out,B6,u53_bout,u55_sout,u54_out,u54_bout,u54_sout);
UnitCell u55(u46_out,1'b0,u54_bout,~u55_bout,u55_out,u55_bout,u55_sout);

assign Q0 = ~u55_bout;

endmodule