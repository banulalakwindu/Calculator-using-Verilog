module non_decoder(output [7:0] dispOut);

//outputs
assign dispOut[0] = 1;
assign dispOut[1] = 1;
assign dispOut[2] = 1;
assign dispOut[3] = 1;
assign dispOut[4] = 1;
assign dispOut[5] = 1;
assign dispOut[6] = 1;
assign dispOut[7] = 1;

endmodule